library ieee;
use ieee.std_logic_1164.all;

library work;
use work.defines.all;

entity map_draws_textures is
	port(
		texture_id : in integer range 0 to 32-1;
		x          : in integer range 0 to 8-1;
		y          : in integer range 0 to 8-1;
		ARGB       : out VGA_ARGB_t
	);
end map_draws_textures;

architecture RTL of map_draws_textures is
	subtype color_t is std_logic_vector(2 downto 0);
	type st is array (0 to 31*8*8-1) of color_t;
	constant c_memory : st := (

		--canto 1 doubleline 0

		"000","000","001","001","001","001","001","001",
		"000","001","000","000","000","000","000","000",
		"001","000","000","000","001","001","001","001",
		"001","000","000","001","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",

		-- canto2 doubleline 1

		"001","001","001","001","001","001","000","000",
		"000","000","000","000","000","000","001","000",
		"001","001","001","001","000","000","000","001",
		"000","000","000","000","001","000","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",

		--canto 3 doubleline 2

		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","000","001","000","000","000","000",
		"001","000","000","000","001","001","001","001",
		"000","001","000","000","000","000","000","000",
		"000","000","001","001","001","001","001","001",

		--canto 4 doubleline 3

		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","001","000","000","001",
		"001","001","001","001","000","000","000","001",
		"000","000","000","000","000","000","001","000",
		"001","001","001","001","001","001","000","000",

		--linha horizont 4

		"001","001","001","001","001","001","001","001",
		"000","000","000","000","000","000","000","000",
		"001","001","001","001","001","001","001","001",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

		-- 5

		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",

		--BLACK-6

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

			--linha horizont 2-*7

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"001","001","001","001","001","001","001","001",
		"000","000","000","000","000","000","000","000",
		"001","001","001","001","001","001","001","001",

		--	linha vert esq  8

		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",

		--margin str8 corner lft 9

		"001","001","001","001","001","001","001","001",
		"000","000","000","000","000","000","000","000",
		"001","001","001","000","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",

		--margin str8 corner rght 10

		"001","001","001","001","001","001","001","001",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","001","001",
		"000","000","000","000","000","001","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",

		-- other vertical 11

		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",

				--map corner1 lft 12

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","001","001",
		"000","000","000","000","000","001","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",

				--map corner2 lft 13

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"001","001","000","000","000","000","000","000",
		"000","000","001","000","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",

				--map corner3 lft 14

		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","001","000","000","000","000","000",
		"001","001","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

				--map corner4 lft 15

		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","001","000","000","000",
		"000","000","000","000","000","001","000","000",
		"000","000","000","000","000","000","001","001",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

		-- str8t single line hori 16

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"001","001","001","001","001","001","001","001",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

		--str8 snglelin vert 17

		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",
		"000","000","000","001","000","000","000","000",

			--ghostbox corner 1 18

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","001","001","001",
		"000","000","000","000","000","001","000","000",
		"000","000","000","000","000","001","000","001",

			--ghost box white 19

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"111","111","111","111","111","111","111","111",
		"111","111","111","111","111","111","111","111",
		"111","111","111","111","111","111","111","111",

					--ghostbox corner 2 20

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"001","001","001","000","000","000","000","000",
		"000","000","001","000","000","000","000","000",
		"001","000","001","000","000","000","000","000",

					--ghostbox corner 3 21

		"000","000","000","000","000","001","000","000",
		"000","000","000","000","000","001","000","000",
		"000","000","000","000","000","001","001","001",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

					--ghostbox corner 4 22

		"000","000","001","000","000","000","000","000",
		"000","000","001","000","000","000","000","000",
		"001","001","001","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

				--map corner1 lft 23

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","001",
		"000","000","000","000","000","000","001","000",
		"000","000","000","000","000","001","000","000",

				--map corner2 lft 24

		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"001","000","000","000","000","000","000","000",
		"000","001","000","000","000","000","000","000",
		"000","000","001","000","000","000","000","000",

				--map corner3 lft 25

		"000","000","001","000","000","000","000","000",
		"000","001","000","000","000","000","000","000",
		"001","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

				--map corner4 lft 26

		"000","000","000","000","000","001","000","000",
		"000","000","000","000","000","000","001","000",
		"000","000","000","000","000","000","000","001",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",
		"000","000","000","000","000","000","000","000",

					--map corner4 lft 27

		"000","001","000","000","000","000","000","000",
		"000","001","000","000","000","000","000","000",
		"000","001","000","000","000","000","000","000",
		"000","001","000","000","000","000","000","000",
		"000","001","000","000","000","001","001","001",
		"000","001","000","000","001","000","000","000",
		"000","001","000","001","000","000","000","000",
		"000","001","000","001","000","000","000","000",

					--map corner4 lft 28

		"000","001","000","001","000","000","000","000",
		"000","001","000","001","000","000","000","000",
		"000","001","000","001","000","000","000","000",
		"000","001","000","000","001","000","000","000",
		"000","001","000","000","000","001","001","001",
		"000","001","000","000","000","000","000","000",
		"000","001","000","000","000","000","000","000",
		"000","001","000","000","000","000","000","000",

					--map corner4 lft 29

		"000","000","000","000","000","000","000","001",
		"000","000","000","000","000","000","000","001",
		"000","000","000","000","000","000","000","001",
		"000","000","000","000","000","000","000","001",
		"001","001","001","001","000","000","000","001",
		"000","000","000","000","001","000","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",

					--map corner4 lft 30

		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","000","001","000","001",
		"000","000","000","000","001","000","000","001",
		"001","001","001","001","000","000","000","001",
		"000","000","000","000","000","000","000","001",
		"000","000","000","000","000","000","000","001",
		"000","000","000","000","000","000","000","001"

	);

begin

	process(texture_id, x, y)
	begin
		if (texture_id = 31) then
			ARGB <= "0000";
		else
			ARGB <= "1" & c_memory((texture_id * 8 * 8 + x + y * 8));
		end if;
	end process;
	
end RTL;
