library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

library work;
use work.defines.all;

entity num_rom is
	port(
		x          :  in integer range 0 to 8-1;
		y          :  in integer range 0 to 8-1;
		texture_id :  in integer range 0 to 10-1;
		ARGB       : out VGA_ARGB_t
	);

end num_rom;

architecture RTL of num_rom is 
signal s_dataout : integer range 0 to 1;
subtype t is integer range 0 to 1;
type st is array (0 to (10*8*8)-1) of t;

constant c_memory : st := 
(
0,1,1,1,1,1,1,0,
0,1,1,1,1,1,1,0,
0,1,0,0,1,1,1,0,
0,1,0,0,1,0,1,0,
0,1,0,1,1,0,1,0,
0,1,1,1,0,0,1,0,
0,1,1,0,0,0,1,0,
0,1,1,1,1,1,1,0,


0,0,0,0,1,0,0,0,
0,0,0,1,1,0,0,0,
0,0,1,1,1,0,0,0,
0,1,1,1,1,0,0,0,
1,1,0,1,1,0,0,0,
0,0,0,1,1,0,0,0,
0,0,0,1,1,0,0,0,
0,1,1,1,1,1,1,0,

0,0,1,1,1,1,0,0,
0,1,1,1,1,1,1,0,
0,1,0,0,0,0,1,0,
0,1,0,0,0,0,1,0,
0,0,0,1,1,1,1,0,
0,1,1,1,1,1,0,0,
0,1,0,0,0,0,0,0,
0,1,1,1,1,1,1,1,


0,1,1,1,1,1,1,0,
0,0,0,0,0,0,0,1,
0,0,0,0,0,0,0,1,
0,1,1,1,1,1,1,0,
0,1,1,1,1,1,1,0,
0,0,0,0,0,0,1,0,
0,0,0,0,0,0,0,1,
0,1,1,1,1,1,1,0,


0,0,0,1,1,1,1,0,
0,0,1,1,1,1,1,0,
0,1,1,0,0,1,1,0,
0,1,0,0,0,1,1,0,
0,1,1,1,1,1,1,0,
0,1,1,1,1,1,1,0,
0,0,0,0,0,1,1,0,
0,0,0,0,0,1,1,0,


0,1,1,1,1,1,1,0,
0,1,1,1,1,1,1,0,
0,1,0,0,0,0,0,0,
0,1,0,0,0,0,0,0,
0,1,1,1,1,1,1,0,
0,0,0,0,0,0,1,0,
0,0,0,0,0,0,1,0,
0,1,1,1,1,1,1,0,


0,0,1,1,1,1,1,0,
0,1,1,0,0,0,1,0,
0,1,0,0,0,0,0,0,
0,1,0,1,1,1,0,0,
0,1,1,1,1,1,1,0,
0,1,0,0,0,0,1,0,
0,1,0,0,0,0,1,0,
0,0,1,1,1,1,0,0,


1,1,1,1,1,1,1,0,
1,1,1,1,1,1,1,0,
0,0,0,0,0,1,1,0,
0,0,0,0,0,1,1,0,
0,0,0,0,0,1,1,0,
0,0,0,0,0,1,1,0,
0,0,0,0,0,1,1,0,
0,0,0,0,0,1,1,0,



0,1,1,1,1,1,1,0,
0,1,0,0,0,0,1,0,
0,1,0,0,0,0,1,0,
0,1,1,1,1,1,1,0,
0,1,1,1,1,1,1,0,
0,1,0,0,0,0,1,0,
0,1,0,0,0,0,1,0,
0,1,1,1,1,1,1,0,

0,1,1,1,1,1,1,0,
0,1,1,1,1,1,1,0,
0,1,0,0,0,0,1,0,
0,1,0,0,0,0,1,0,
0,1,1,1,1,1,1,0,
0,0,0,0,0,0,1,0,
0,0,0,0,0,0,1,0,
0,1,1,1,1,1,1,0

);

begin

	s_dataout <= c_memory(texture_id * 8 * 8 + x + y * 8);

	color_map : process(s_dataout)
	begin
		if (s_dataout = 1) then
			ARGB <= "1111";
		else
			ARGB <= "0000";
		end if ;
	end process;

end;